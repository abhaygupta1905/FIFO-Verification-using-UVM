import uvm_pkg::*; 
 
`include "seq_item.sv" 
`include "base_seq.sv" 
`include "sequencer.sv" 
`include "driver.sv" 
`include "monitor.sv" 
`include "scoreboard.sv" 
`include "agent.sv" 
`include "env.sv" 
`include "base_test.sv"
